dut_top
